interface intf(input logic clk,resetn);
  
  //declaring the signals
  logic Rqst0;
  logic Rqst1;
  logic Rqst2;
  logic Rqst3;
logic Grant0;
  logic Grant1;
  logic Grant2;
  logic Grant3;

  
endinterface
